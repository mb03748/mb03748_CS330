module tb2
(


);
