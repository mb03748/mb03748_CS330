module top
  (
  
  ):
  
  wire a;
  wire b;
  wire CarryIn;
  wire [3:0]ALUop;
  reg Result;
  reg CarryOut;
  